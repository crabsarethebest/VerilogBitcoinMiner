module hello_world ();

logic x = 1'b1;
endmodule
